LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY override_controller IS
	-- CONSTANTES
	GENERIC (
		CONSTANT OPERATION_DISTANCE : INTEGER := 136; --140 1; -- Minimum aantal PWM pulsen die gepasseerd moeten zijn sinds het uitvoeren van de vorige mogelijkheid van de override controller
		CONSTANT FORWARD_PWM_COUNT : INTEGER := 20;--20; -- Aantal PWM pulsen dat die in de staten forward, left, en right moet doorbrengen
		CONSTANT LEFT_PWM_COUNT : INTEGER := 40;--35;
		CONSTANT RIGHT_PWM_COUNT : INTEGER := 55; --35;
		CONSTANT TX_MIJN : std_logic_vector(7 DOWNTO 0) := "00110000";
		CONSTANT TX_GEEN_MIJN : std_logic_vector(7 DOWNTO 0) := "00110001";
		CONSTANT RELATIVE_SEND : INTEGER := 20;--20;
		CONSTANT DISTANCE_ON_RESET : unsigned := "00000010010110";-- waarde van de distance_counter na een systeemreset
		CONSTANT MINE_FORWARD : INTEGER := 12
	);

	PORT (
		clk, reset            : IN std_logic;
		translator_out        : IN std_logic_vector(7 DOWNTO 0);
		override_vector       : OUT std_logic_vector(3 DOWNTO 0);
		override              : OUT std_logic;
		translator_out_reset  : OUT std_logic;
		count_reset           : IN std_logic;
		sensor_l              : IN std_logic;
		sensor_m              : IN std_logic;
		sensor_r              : IN std_logic;
		tx_out                : OUT std_logic_vector(7 DOWNTO 0);
		tx_send_out           : OUT std_logic;
		count_in              : IN std_logic_vector (19 DOWNTO 0);
 
		an                    : OUT STD_LOGIC_VECTOR (3 DOWNTO 0); -- Selectie van schermpje
		sseg                  : OUT STD_LOGIC_VECTOR (7 DOWNTO 0); -- Getal dat weergegeven moet worden.
		led                   : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		mine_button           : IN std_logic
	);
END ENTITY override_controller;

ARCHITECTURE behavioural OF override_controller IS
	-- TYPES
	TYPE override_controller_states IS (-- Mogelijkheden override controller
	read_sensor_and_listen, 
	forward, 
	right90, right, fastright, 
	left90, left, fastleft, 
	forward_station, left_station, right_station, mine);
	TYPE station_state_type IS (-- Staten binnen een opdracht zoals een bocht naar links of een station aan de voorkant.
	first2, first, second, third, fourth, fifth);
	TYPE tx_state IS (-- Staten gebruikt bij de transmitter
	tx_idle, tx_wait_normal, tx_send);

	TYPE prev_directiontype IS(left, right, forward);

	-- Controle var
 
	SIGNAL prev_direction, next_prev_direction : prev_directiontype; --Om de vorige richting bij te houden. Is nodig voor een efficiente de bocht na een detectie van een mijn.
	SIGNAL station_state, new_station_state : station_state_type; 
	SIGNAL override_cont_state, override_cont_new_state : override_controller_states; 
	SIGNAL tx_state_reg, tx_state_next : tx_state; 
	SIGNAL pwm_count, new_pwm_count, distance_count, new_distance_count : unsigned (13 DOWNTO 0); -- Geheugenelementen voor de pwm-tellers voor de bochten en voor de afstand lijnengevolgd
	SIGNAL pwm_count_out : std_logic_vector (13 DOWNTO 0);
	SIGNAL pwm_count_reset, distance_count_reset : std_logic; -- Resets voor de pwm-tellers.
	SIGNAL next_translator_out_reset : std_logic;
 
	--signalen voor display
	SIGNAL override_state_sseg, station_state_sseg : STD_LOGIC_VECTOR (7 DOWNTO 0);
 
BEGIN
PROCESS (clk, reset) -- Check op rising edge en op resets
BEGIN
	IF (rising_edge(clk)) THEN
		IF (reset = '1') THEN
			override_cont_state <= read_sensor_and_listen; -- Zet de states in de eerste staat
			station_state <= first;
			tx_state_reg <= tx_idle;
			translator_out_reset <= '0';
			prev_direction <= forward;
		ELSE
			override_cont_state <= override_cont_new_state; -- Ga naar de volgende staat op de rising edge
			station_state <= new_station_state;
			tx_state_reg <= tx_state_next;
			translator_out_reset <= next_translator_out_reset;
			prev_direction <= next_prev_direction;
		END IF;
	END IF;
END PROCESS;

PROCESS (clk, translator_out, sensor_l, sensor_m, sensor_r, override_cont_state, pwm_count, distance_count, pwm_count_out, station_state, prev_direction, mine_button) -- Gedrag van specefieke handelingen
BEGIN
	next_prev_direction <= prev_direction;
	next_translator_out_reset <= '0';
	new_station_state <= station_state;
	pwm_count_reset <= '0';
	CASE override_cont_state IS
		WHEN read_sensor_and_listen => -- In deze staat zal hij lijnvolgen (dwz, overide = 0) totdat een bepaalde afstand is overschreden
			-- EN de sensoren allemaal zwart zijn (Bij een kruispunt!)
 
			distance_count_reset <= '0'; -- De distance-teller telt gewoon door
			override_vector <= "0000"; -- Stel hij override de controller hier, dan zet hij de robot stil.
			new_station_state <= first; -- Eerste staat in de station FSM, (als het ware een reset van deze FSM)
 
 

			IF (sensor_l = '0' AND sensor_m = '0' AND sensor_r = '0' AND distance_count > OPERATION_DISTANCE) THEN -- neem de lijnvolger over.
				override <= '1'; 
 
				next_translator_out_reset <= '1';
				pwm_count_reset <= '1'; -- Hij komt in de override stand en mag beginnen met tellen van het aantal pwm perioden. Deze teller is voor de bochten.
				CASE translator_out IS -- Afhankelijk van het ingekomen signaal van C wordt er hier gekozen uit de juiste bocht.
					WHEN "10000001" => override_cont_new_state <= forward;
					WHEN "10000010" => override_cont_new_state <= right;
					WHEN "10000100" => override_cont_new_state <= left;
					WHEN "11000001" => override_cont_new_state <= forward_station;
					WHEN "11000010" => override_cont_new_state <= right_station;
					WHEN "11000100" => override_cont_new_state <= left_station;
					WHEN OTHERS => override_cont_new_state <= read_sensor_and_listen;
						next_translator_out_reset <= '0'; --Voor als er nog geen nieuwe opdracht binnen is (translator_out = "00000000"). Dan geen translator_out_reset doen en blijven wachten.
				END CASE;
			ELSE
				override <= '0';
				pwm_count_reset <= '0'; -- pwm_count is een counter die telt per 20 ms. Zo is het aantal pwm pulsen te tellen.
				override_cont_new_state <= read_sensor_and_listen;
			END IF;
 
			IF (Mine_button = '1') THEN --als een mijn gevonden is naar de mijn staat gaan.
				pwm_count_reset <= '1';
				override <= '1';
				override_cont_new_state <= mine;
				next_translator_out_reset <= '1';
			END IF;

			-- Dit zijn de staten voor de verschillende bochten: rechtdoor, links en rechts bij een kruising.
			-- Er zijn ook staten voor een bocht naar een station, hier zal de staat ook de bocht aan het einde van de weg maken.
			-- Ook de mijn staat staat hier bij.
			-- Aan het einde van de actie komt de override_controller weer in zijn read_sensor_and_listen staat.

		WHEN forward => --Een korte periode vooruit rijden en daarna weer over op lijnvolgen.
			next_prev_direction <= forward;
			CASE station_state IS 
				WHEN first => 
					distance_count_reset <= '0'; -- Reset de beide tellers niet
					pwm_count_reset <= '0';
					override <= '0'; -- Gewoon lijnvolgen, hij zal automatisch recht door rijden!
					override_vector <= "0001"; -- vooruit
					override_cont_new_state <= forward; -- blijf in forward
 
					IF (unsigned(pwm_count_out) < FORWARD_PWM_COUNT) THEN -- Zie lijst met constantes
						new_station_state <= first; -- Blijf in dezelfde staat als hij nog niet lang genoeg rechtdoor heeft gereden
					ELSE
						new_station_state <= second; -- Ga naar de volgende staat
					END IF;
				WHEN OTHERS => --second and others.
					distance_count_reset <= '1'; -- Reset de gereden afstand staat
					pwm_count_reset <= '1'; -- Reset de counter voor de handelingen
					override <= '0'; -- Lijnvolgen
					override_vector <= "0000";-- Moet iets zijn, dont care
					override_cont_new_state <= read_sensor_and_listen; -- Ga naar de begin staat

			END CASE;
 
		WHEN left => -- Voor een bepaalde tijd een bocht naar links maken en daarna weer lijnvolgen.
			next_prev_direction <= left;
			distance_count_reset <= '0';
			pwm_count_reset <= '0'; 
			override_cont_new_state <= left;
			override_vector <= "0000";

			CASE station_state IS
			
								WHEN first =>
					override <= '0';
					IF (unsigned(pwm_count_out) < 14) THEN -- Zie lijst met constantes
						new_station_state <= first; -- Blijf in dezelfde staat als hij nog niet lang genoeg rechtdoor heeft gereden
					ELSE
						new_station_state <= first2; -- Ga naar de volgende staat
					END IF;
					
					
				WHEN first2 => 
					override <= '1';
					override_vector <= "0111"; -- harde bocht naar links 0111
					IF (unsigned(pwm_count_out) < LEFT_PWM_COUNT) THEN
						new_station_state <= first2; -- Blijf in dezelfde staat
					ELSE
						new_station_state <= second; -- Ga naar de volgende
					END IF;
				WHEN second => -- Rechtdoor rijden tot dat de linker sensor weer de lijn ziet. Dit geeft de soepelste bocht.
					override <= '1';
					override_vector <= "0001"; -- rechtdoor

					IF (sensor_l = '0') THEN 
						new_station_state <= third; -- ga naar volgende staat
					ELSE
						new_station_state <= second; --blijf in dezelfde staat
					END IF;
 
				WHEN OTHERS => --second and others.
					distance_count_reset <= '1'; -- Reset de gereden distance, deze is zo weer nodig
					pwm_count_reset <= '1'; -- Reset de handelings pwm-teller
					override <= '0'; -- Lijnvolen
					override_vector <= "0000";
					override_cont_new_state <= read_sensor_and_listen;

			END CASE;
			
			IF (Mine_button = '1') THEN --als een mijn gevonden is naar de mijn staat gaan.
				pwm_count_reset <= '1';
				override <= '1';
				override_cont_new_state <= mine;
				next_translator_out_reset <= '1';
			END IF;
			
		WHEN right => -- Voor een bepaalde periode een bocht naar rechts maken en dan weer lijnvolgen.
			next_prev_direction <= right;
			distance_count_reset <= '0';
			pwm_count_reset <= '0';
			override_cont_new_state <= right;
			override_vector <= "0000";

			CASE station_state IS
			
					WHEN first =>
					override <= '0';
					IF (unsigned(pwm_count_out) < 14) THEN -- Zie lijst met constantes
						new_station_state <= first; -- Blijf in dezelfde staat als hij nog niet lang genoeg rechtdoor heeft gereden
					ELSE
						new_station_state <= first2; -- Ga naar de volgende staat
					END IF;
					
				WHEN first2 => 
					override <= '1';
					override_vector <= "0100"; -- harde bocht naar rechts

					IF (unsigned(pwm_count_out) < RIGHT_PWM_COUNT) THEN
						new_station_state <= first2;
					ELSE
						new_station_state <= second;
					END IF;
 
				WHEN second => -- Rechtdoor rijden tot dat de rechter sensor weer de lijn ziet. Dit geeft de soepelste bocht.
					override <= '1';
					override_vector <= "0001"; -- rechtdoor
					IF (sensor_r = '0') THEN -- oud: NOT(sensor_l = '0' AND sensor_m = '0')
						new_station_state <= third;
					ELSE
						new_station_state <= second;
					END IF; 
 
				WHEN OTHERS => --second and others.
					distance_count_reset <= '1';
					pwm_count_reset <= '1';
					override <= '0';
					override_vector <= "0000";
					override_cont_new_state <= read_sensor_and_listen;
 
			END CASE;
			
		IF (Mine_button = '1') THEN --als een mijn gevonden is naar de mijn staat gaan.
				pwm_count_reset <= '1';
				override <= '1';
				override_cont_new_state <= mine;
				next_translator_out_reset <= '1';
			END IF; 
	
		WHEN left_station => 
			distance_count_reset <= '0';
			pwm_count_reset <= '0';
			override_vector <= "1000";
			override_cont_new_state <= left_station;
			override_cont_new_state <= left_station;
			CASE station_state IS
				WHEN first => -- Gewoon de bocht naar links(gekopierd)
					
					override <= '1';
					override_vector <= "0111"; -- harde bocht naar links
 
					IF (unsigned(pwm_count_out) < LEFT_PWM_COUNT) THEN
						new_station_state <= first;
					ELSE
						new_station_state <= second;
					END IF;
				WHEN second => -- De lijn terugvinden door rechtdoor te rijden.
					override <= '1';
					override_vector <= "0001"; -- Rechtdoor
 
					IF (sensor_r = '0' AND sensor_m = '0') THEN
						new_station_state <= THIRD;
					ELSE
						new_station_state <= second;
					END IF;
 
				WHEN third => --lijnvolgen (override = '0') zolang in ieder geval 1 van de sensoren een lijn ziet. Zo rijd hij tot het einde van de lijn (waar ze alle drie wit (='1') worden)
					override <= '0';
					IF (sensor_l = '0' OR sensor_m = '0' OR sensor_r = '0') THEN
						new_station_state <= third;
					ELSE
						new_station_state <= fourth;
					END IF;
				WHEN fourth => --Bocht maken als hij aan het einde van de lijn is. Dan geldt: sensor_l ='1' (wit). Dan 180 graden RECHTSOM draaien. De linker sensor zal als laatste weer zwart worden. Dan verder naar de volgende stap.
					override <= '1';
					override_vector <= "0100"; -- drive_motor_fastright.
					IF (sensor_l = '1') THEN
						new_station_state <= fourth;
					ELSE
						new_station_state <= fifth;
					END IF;
				WHEN fifth => -- De robot is klaar om weer lijn te volgen, hij verlaat de override stand.
					distance_count_reset <= '0'; -- In het geval dat de robot een station bezocht heeft hoeft hij niet de distance counter te resetten, omdat hij geen zwarte stip meer tegen zal komen.
					pwm_count_reset <= '1';
					override <= '0';
					override_cont_new_state <= read_sensor_and_listen;
					new_station_state <= first;
					
					
					
					WHEN OTHERS => 
										distance_count_reset <= '0'; -- In het geval dat de robot een station bezocht heeft hoeft hij niet de distance counter te resetten, omdat hij geen zwarte stip meer tegen zal komen.
					pwm_count_reset <= '1';
					override <= '0';
					override_cont_new_state <= read_sensor_and_listen;
					new_station_state <= first;
					
			END CASE;

		WHEN forward_station => 
			distance_count_reset <= '0';
			pwm_count_reset <= '0';
			override_vector <= "1000"; 
			override_cont_new_state <= forward_station;
			CASE station_state IS
				WHEN first => -- Lijnvolgen
					override <= '0';
					IF (sensor_l = '0' OR sensor_m = '0' OR sensor_r = '0') THEN --lijnvolgen zolang in ieder geval 1 van de sensoren een lijn ziet. Zo rijd hij tot het einde van de lijn (waar ze alle drie wit (='1') worden)
						new_station_state <= first;
					ELSE
						new_station_state <= second;
					END IF;
				WHEN second => --Bocht maken als hij aan het einde van de lijn is. Dan geldt: sensor_l ='1' (wit). Dan 180 graden RECHTSOM draaien. De linker sensor zal als laatste weer zwart worden. Dan verder naar de volgende stap.
					override <= '1';
					override_vector <= "0100"; -- drive_motor_right90.
					IF (sensor_l = '1') THEN
						new_station_state <= second;
					ELSE
						new_station_state <= third;
					END IF;
				WHEN others => -- De robot is klaar om weer lijn te volgen, hij verlaat de override stand. Hij moet hier weer een signaal sturen naar de pc dat hij het volgende commando wil.
					pwm_count_reset <= '1';
					override <= '0';
					override_cont_new_state <= read_sensor_and_listen;
					new_station_state <= first;
			END CASE;

		WHEN right_station => 
			distance_count_reset <= '0';
			pwm_count_reset <= '0';
			override_vector <= "1000";
			override_cont_new_state <= right_station;
			CASE station_state IS
				WHEN first => -- Gewoon de bocht naar rechts (gekopierd)
					override <= '1';
					override_vector <= "0100"; -- harde bocht naar links
 
					IF (unsigned(pwm_count_out) < RIGHT_PWM_COUNT) THEN
						new_station_state <= first;
					ELSE
						new_station_state <= second;
					END IF;
				WHEN second => 
					override <= '1';
					override_vector <= "0001"; -- Vooruit om de lijn terug te vinden.
					IF (sensor_l = '0' AND sensor_m = '0') THEN
						new_station_state <= THIRD;
					ELSE
						new_station_state <= second;
					END IF;
 
				WHEN third => --lijnvolgen (override = '0') zolang in ieder geval 1 van de sensoren een lijn ziet. Zo rijd hij tot het einde van de lijn (waar ze alle drie wit (='1') worden)
					override <= '0';
					IF (sensor_l = '0' OR sensor_m = '0' OR sensor_r = '0') THEN
						new_station_state <= third;
					ELSE
						new_station_state <= fourth;
					END IF;
				WHEN fourth => --Bocht maken als hij aan het einde van de lijn is. Dan geldt: sensor_l ='1' (wit). Dan 180 graden LINKSOM draaien. De linker sensor zal als laatste weer zwart worden. Dan verder naar de volgende stap.
					override <= '1';
					override_vector <= "0111"; -- drive_motor_left90.
					IF (sensor_r = '1') THEN
						new_station_state <= fourth;
					ELSE
						new_station_state <= fifth;
					END IF;
				WHEN fifth => -- De robot is klaar om weer lijn te volgen, hij verlaat de override stand.
					distance_count_reset <= '0'; -- In het geval dat de robot een station bezocht heeft hoeft hij niet de distance counter te resetten, omdat hij geen zwarte stip meer tegen zal komen.
					pwm_count_reset <= '1';
					override <= '0';
					override_cont_new_state <= read_sensor_and_listen;
					new_station_state <= first;
					
					WHEN OTHERS => 
										distance_count_reset <= '0'; -- In het geval dat de robot een station bezocht heeft hoeft hij niet de distance counter te resetten, omdat hij geen zwarte stip meer tegen zal komen.
					pwm_count_reset <= '1';
					override <= '0';
					override_cont_new_state <= read_sensor_and_listen;
					new_station_state <= first;
			END CASE;
 
		WHEN mine => 
			distance_count_reset <= '0';
			pwm_count_reset <= '0';
			override_vector <= "1000"; -- moet iets zijn
			override_cont_new_state <= mine;
			CASE station_state IS
			
				WHEN  first => --Klein stukje nog lijnvolgen.
					override <= '0';
					IF (unsigned(pwm_count_out) < MINE_FORWARD) THEN
						new_station_state <= first;
					ELSE
						new_station_state <= second;
					END IF;
				
				WHEN second =>  --Om de as draaien. Afhankelijk van de vorige richting dit linksom of rechtsom doen
					override <= '1';
					IF (prev_direction = forward) THEN
						override_vector <= "0100"; --right90
					ELSIF (prev_direction = right) THEN--OM!!!
						override_vector <= "0111"; --left90
					ELSE --prev = left
						override_vector <= "0100"; --right90
					END IF;
 
					IF (unsigned(pwm_count_out) < 90) THEN -- om as draaien zolang tenminste een van de sensoren de lijn nog ziet. Daarna word alles wit en gaat hij naar de volgende staat.
						new_station_state <= second;
					ELSE
						new_station_state <= third;
					END IF;
 
 
				WHEN third => -- Om as draaien in zelfde richting als in staat 'second'. Nu door draaien tot de sensoren weer de lijn zien.
					override <= '1';
					IF (prev_direction = forward) THEN
						override_vector <= "0100"; --right90
						IF (sensor_r = '0') THEN
							new_station_state <= fourth; 
						ELSE
							new_station_state <= third;
						END IF;
					ELSIF (prev_direction = right) THEN --OM!!!
						override_vector <= "0111"; -- left90
						IF (sensor_l = '0') THEN
							new_station_state <= fourth; 
						ELSE
							new_station_state <= third;
						END IF;
					ELSE --prev = left
						override_vector <= "0100"; -- right90
						IF (sensor_r = '0') THEN --OM!!!
							new_station_state <= fourth;
						ELSE
							new_station_state <= third;
						END IF;
					END IF;
 
				WHEN OTHERS => --lijn is teruggevonden en override controller kan terug naar read_sensor_and_listen staat.
					override <= '0';
					distance_count_reset <= '0';
					pwm_count_reset <= '1';
					override_cont_new_state <= read_sensor_and_listen;
 
					new_station_state <= first;
 
 
			END CASE;

		WHEN OTHERS => 
			distance_count_reset <= '0';
			pwm_count_reset <= '0';
			override <= '0';
			override_vector <= "0000";-- moet iets zijn
			override_cont_new_state <= read_sensor_and_listen;

	END CASE;
END PROCESS;

-- Counter van PWM perioden (20 ms). Wordt gebruikt voor bochten van een bepaalde lengte
PROCESS (count_reset, pwm_count_reset, reset, clk)
BEGIN
	IF (reset = '1' OR pwm_count_reset = '1') THEN
		pwm_count <= (OTHERS => '0');
	ELSIF (rising_edge(count_reset)) THEN
		pwm_count <= new_pwm_count;
	END IF;
END PROCESS;

PROCESS (pwm_count)
BEGIN
	new_pwm_count <= pwm_count + 1;
END PROCESS;
pwm_count_out <= std_logic_vector(pwm_count);

-- Counter van PWM perioden, maar dan voor de afstandsmeting (Het stukje tussen de twee stations)
PROCESS (count_reset, distance_count_reset, reset, clk)
BEGIN
	IF (reset = '1') THEN
		distance_count <= DISTANCE_ON_RESET; -- Bij een reset doet de distance counter er niet toe, hij begint dan namelijk bij een station.
	ELSIF (distance_count_reset = '1') THEN
		distance_count <= (OTHERS => '0');
	ELSIF (rising_edge(count_reset)) THEN
		distance_count <= new_distance_count;
	END IF;
END PROCESS;

PROCESS (distance_count)
BEGIN
	new_distance_count <= distance_count + 1;
END PROCESS;

-- tx signalen. Zal versturen op het kruisen van de stip tussen de kruispunten, of bij het verschijnen in een *_station staat
PROCESS (clk, sensor_l, sensor_r, sensor_m, distance_count, distance_count_reset, override_cont_state, tx_state_reg, mine_button)
BEGIN
	tx_state_next <= tx_state_reg;
	tx_out <= TX_GEEN_MIJN;
 
	IF (mine_button = '1' and tx_state_reg /= tx_wait_normal) THEN
		tx_out <= TX_MIJN;
		tx_state_next <= tx_send;
	END IF;
 
	CASE(tx_state_reg) IS
	WHEN tx_idle => -- Wachten wachten wachten wachten....
	tx_send_out <= '0';
	IF (override_cont_state /= read_sensor_and_listen) THEN
		tx_state_next <= tx_send;
	END IF;
	WHEN tx_send => -- stuur 1 klokpuls
	tx_send_out <= '1';
	tx_state_next <= tx_wait_normal;
 
	WHEN tx_wait_normal => -- Forceer hem om maar een keer te sturen bij normale states. Aan het einde van een handeling wordt distance_count gereset
	tx_send_out <= '0';
	IF (override_cont_state = read_sensor_and_listen) THEN
		tx_state_next <= tx_idle;
	END IF;
END CASE;
END PROCESS;


--Segmentendisplay aansturen
PROCESS (station_state_sseg, override_state_sseg, distance_count, count_in) --Multiplexer. Zet om en om een waarde op een van de displays.
BEGIN
sseg(7) <= '0'; --decimale punt uit
IF (count_in(15) = '0') THEN --Count_in, de teller van de 50Mhz clock, word gebruikt om te multiplexen. De frequentie is: (50*10^6)/(2^15) = 1526 Hz
	an <= "1110";
	sseg <= override_state_sseg;
ELSE
	sseg <= station_state_sseg;
	an <= "0111";
END IF;
END PROCESS;

WITH translator_out SELECT
override_state_sseg(7 DOWNTO 0) <= 
	"01000000" WHEN "00000000", --0 leeg
	"01111001" WHEN "10000001", --1 vooruit
	"00100100" WHEN "10000100", --2 links
	"00110000" WHEN "10000010", --3 rechts
	"00011001" WHEN "11000001", --4 voorruit station
	"00010010" WHEN "11000100", --5 links station
	"00000010" WHEN "11000010", --6 rechts station
	"01111000" WHEN "10000000", --7 stop
	"00001110" WHEN OTHERS; --f
 
WITH station_state SELECT
station_state_sseg(7 DOWNTO 0) <= 
	"01111001" WHEN first, --1
	"00100100" WHEN second, --2
	"00110000" WHEN third, --3
	"00011001" WHEN fourth, --4
	"00010010" WHEN fifth, --5
	"00001110" WHEN OTHERS; --f

 
--Leds aansturen
PROCESS (distance_count)
BEGIN
IF (distance_count < 18) THEN --18
	led <= "00000000";
ELSIF (distance_count < 36) THEN -- 36
	led <= "00000001";
ELSIF (distance_count < 54) THEN -- 54
	led <= "00000011";
ELSIF (distance_count < 72) THEN -- 72
	led <= "00000111";
ELSIF (distance_count < 90) THEN -- 90
	led <= "00001111";
ELSIF (distance_count < 108) THEN --108
	led <= "00011111";
ELSIF (distance_count < 126) THEN --126
	led <= "00111111"; 
ELSIF (distance_count < operation_distance) THEN -- 144
	led <= "01111111";
ELSE
	led <= "11111111";
END IF;

END PROCESS;
END ARCHITECTURE behavioural;